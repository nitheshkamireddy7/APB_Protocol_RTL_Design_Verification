module APB_master (

  
);
endmodule
